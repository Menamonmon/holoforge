module cocotb_iverilog_dump();
initial begin
    $dumpfile("/Users/yabi/Documents/Schooly_Stuff/6.111/holoforge/sim/sim_build/mig_write_req_generator.fst");
    $dumpvars(0, mig_write_req_generator);
end
endmodule
