typedef logic signed [15:0] vfixed_t;
typedef vfixed_t vertex_t[3];
typedef vfixed_t normal_t[3];
typedef logic [7:0] color_id_t;
typedef color_id_t vcolor_t[3];

